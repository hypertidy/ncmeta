netcdf avhrr-only-v2.19810901 {
dimensions:
	time = 1 ;
	zlev = 1 ;
	lat = 10 ;
	lon = 14 ;
variables:
	float time(time) ;
		time:long_name = "Center time of the day" ;
		time:units = "days since 1978-01-01 00:00:00" ;
	float zlev(zlev) ;
		zlev:long_name = "Sea surface height" ;
		zlev:units = "meters" ;
		zlev:actual_range = "0, 0" ;
	float lat(lat) ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:grids = "Uniform grid from -89.875 to 89.875 by 0.25" ;
	float lon(lon) ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:grids = "Uniform grid from 0.125 to 359.875 by 0.25" ;
	short sst(time, zlev, lat, lon) ;
		sst:long_name = "Daily sea surface temperature" ;
		sst:units = "degrees C" ;
		sst:_FillValue = -999s ;
		sst:add_offset = 0.f ;
		sst:scale_factor = 0.01f ;
		sst:valid_min = -300s ;
		sst:valid_max = 4500s ;
	short anom(time, zlev, lat, lon) ;
		anom:long_name = "Daily sea surface temperature anomalies" ;
		anom:units = "degrees C" ;
		anom:_FillValue = -999s ;
		anom:add_offset = 0.f ;
		anom:scale_factor = 0.01f ;
		anom:valid_min = -1200s ;
		anom:valid_max = 1200s ;
	short err(time, zlev, lat, lon) ;
		err:long_name = "Estimated error standard deviation of analysed_sst" ;
		err:units = "degrees C" ;
		err:_FillValue = -999s ;
		err:add_offset = 0.f ;
		err:scale_factor = 0.01f ;
		err:valid_min = 0s ;
		err:valid_max = 1000s ;
	short ice(time, zlev, lat, lon) ;
		ice:long_name = "Sea ice concentration" ;
		ice:units = "percentage" ;
		ice:_FillValue = -999s ;
		ice:add_offset = 0.f ;
		ice:scale_factor = 0.01f ;
		ice:valid_min = 0s ;
		ice:valid_max = 100s ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:title = "Daily-OI-V2, final, Data (Ship, Buoy, AVHRR, GSFC-ice)" ;
		:History = "Version 2.0" ;
		:creation_date = "2011-05-04" ;
		:Source = "NOAA/National Climatic Data Center" ;
		:Contact = "Dick Reynolds, email: Richard.W.Reynolds@noaa.gov & Chunying Liu, email: Chunying.liu@noaa.gov" ;
}
