netcdf pr_2019 {
dimensions:
	lon = 1 ;
	lat = 1 ;
	day = 1 ;
	crs = 1 ;
variables:
	double lon(lon) ;
		lon:units = "degrees_east" ;
		lon:description = "longitude" ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:axis = "X" ;
	double lat(lat) ;
		lat:units = "degrees_north" ;
		lat:description = "latitude" ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:axis = "Y" ;
	double day(day) ;
		day:description = "days since 1900-01-01" ;
		day:units = "days since 1900-01-01 00:00:00" ;
		day:long_name = "time" ;
		day:standard_name = "time" ;
		day:calendar = "gregorian" ;
	ushort crs(crs) ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:long_name = "WGS 84" ;
		crs:inverse_flattening = 298.257223563 ;
		crs:GeoTransform = "-124.7666666333333 0.041666666666666 0  49.400000000000000 -0.041666666666666" ;
		crs:spatial_ref = "GEOGCS[\"WGS 84\",DATUM[\"WGS_1984\",SPHEROID[\"WGS 84\",6378137,298.257223563,AUTHORITY[\"EPSG\",\"7030\"]],AUTHORITY[\"EPSG\",\"6326\"]],PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]],AUTHORITY[\"EPSG\",\"4326\"]]" ;
		crs:_Storage = "chunked" ;
		crs:_ChunkSizes = 1 ;
		crs:_DeflateLevel = 9 ;
		crs:_Endianness = "little" ;
	ushort precipitation_amount(day, lat, lon) ;
		precipitation_amount:_FillValue = 32767US ;
		precipitation_amount:units = "mm" ;
		precipitation_amount:description = "Daily Accumulated Precipitation" ;
		precipitation_amount:long_name = "pr" ;
		precipitation_amount:standard_name = "pr" ;
		precipitation_amount:missing_value = 32767s ;
		precipitation_amount:dimensions = "lon lat time" ;
		precipitation_amount:grid_mapping = "crs" ;
		precipitation_amount:coordinate_system = "WGS84,EPSG:4326" ;
		precipitation_amount:scale_factor = 0.1 ;
		precipitation_amount:add_offset = 0. ;
		precipitation_amount:coordinates = "lon lat" ;
		precipitation_amount:_Unsigned = "true" ;

// global attributes:
		:geospatial_bounds_crs = "EPSG:4326" ;
		:Conventions = "CF-1.6" ;
		:geospatial_bounds = "POLYGON((-124.7666666333333 49.400000000000000, -124.7666666333333 25.066666666666666, -67.058333300000015 25.066666666666666, -67.058333300000015 49.400000000000000, -124.7666666333333 49.400000000000000))" ;
		:geospatial_lat_min = "25.066666666666666" ;
		:geospatial_lat_max = "49.40000000000000" ;
		:geospatial_lon_min = "-124.7666666333333" ;
		:geospatial_lon_max = "-67.058333300000015" ;
		:geospatial_lon_resolution = "0.041666666666666" ;
		:geospatial_lat_resolution = "0.041666666666666" ;
		:geospatial_lat_units = "decimal_degrees north" ;
		:geospatial_lon_units = "decimal_degrees east" ;
		:coordinate_system = "EPSG:4326" ;
		:author = "John Abatzoglou - University of Idaho, jabatzoglou@uidaho.edu" ;
		:date = "01 August 2019" ;
		:note1 = "The projection information for this file is: GCS WGS 1984." ;
		:note2 = "Citation: Abatzoglou, J.T., 2013, Development of gridded surface meteorological data for ecological applications and modeling, International Journal of Climatology, DOI: 10.1002/joc.3413" ;
		:last_permanent_slice = "152" ;
		:last_early_slice = "212" ;
		:last_provisional_slice = "206" ;
		:note3 = "Data in slices after last_permanent_slice (1-based) are considered provisional and subject to change with subsequent updates" ;
		:note4 = "Data in slices after last_provisional_slice (1-based) are considered early and subject to change with subsequent updates" ;
		:note5 = "Days correspond approximately to calendar days ending at midnight, Mountain Standard Time (7 UTC the next calendar day)" ;
		:_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.5" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
}
