netcdf example3 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	X = 1 ;
	Y = 1 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1900-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	float lon(Y, X) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude coordinate" ;
		lon:units = "degrees_east" ;
		lon:_CoordinateAxisType = "Lon" ;
	float lat(Y, X) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude coordinate" ;
		lat:units = "degrees_north" ;
		lat:_CoordinateAxisType = "Lat" ;
	double X(X) ;
		X:standard_name = "projection_x_coordinate" ;
		X:long_name = "x coordinate of projection" ;
		X:units = "meters" ;
		X:axis = "X" ;
	double Y(Y) ;
		Y:standard_name = "projection_y_coordinate" ;
		Y:long_name = "y coordinate of projection" ;
		Y:units = "meters" ;
		Y:axis = "Y" ;
	int ETRS89-LAEA ;
		ETRS89-LAEA:missing_value = -1. ;
		ETRS89-LAEA:grid_mapping_name = "lambert_azimuthal_equal_area" ;
		ETRS89-LAEA:longitude_of_projection_origin = 10. ;
		ETRS89-LAEA:latitude_of_projection_origin = 52. ;
		ETRS89-LAEA:false_easting = 4321000. ;
		ETRS89-LAEA:false_northing = 3210000. ;
		ETRS89-LAEA:inverse_flattening = 298.257222101 ;
		ETRS89-LAEA:semi_major_axis = 6378137. ;
	float pr(time, Y, X) ;
		pr:long_name = "PRECIPITATION" ;
		pr:units = "mm.d-1" ;
		pr:grid_mapping = "ETRS89-LAEA" ;
		pr:coordinates = "lat lon" ;
		pr:_FillValue = -999.99f ;
		pr:missing_value = -999.99f ;
		pr:grid_name = "al05.etrs.laea" ;
		pr:version = "v1.2" ;
		pr:prod_date = "2013-07-15" ;

// global attributes:
		:CDI = "Climate Data Interface version 1.9.1 (http://mpimet.mpg.de/cdi)" ;
		:history = "Thu Oct 04 14:37:21 2018: cdo -C seltimestep,1 /home/esp-shared-a/Observations/EURO4M-APGD/EURO4M-APGD-1971-2008.nc example3.nc\n",
			"Fri Nov  1 13:32:07 2013: ncrename -v PRECIPITATION,pr EURO4M-APGD-1971-2008.nc\n",
			"Fri Nov  1 13:29:54 2013: ncrcat RapdD_al05.etrs.laea_19710100.nc RapdD_al05.etrs.laea_19710200.nc RapdD_al05.etrs.laea_19710300.nc RapdD_al05.etrs.laea_19710400.nc RapdD_al05.etrs.laea_19710500.nc RapdD_al05.etrs.laea_19710600.nc RapdD_al05.etrs.laea_19710700.nc RapdD_al05.etrs.laea_19710800.nc RapdD_al05.etrs.laea_19710900.nc RapdD_al05.etrs.laea_19711000.nc RapdD_al05.etrs.laea_19711100.nc RapdD_al05.etrs.laea_19711200.nc RapdD_al05.etrs.laea_19720100.nc RapdD_al05.etrs.laea_19720200.nc RapdD_al05.etrs.laea_19720300.nc RapdD_al05.etrs.laea_19720400.nc RapdD_al05.etrs.laea_19720500.nc RapdD_al05.etrs.laea_19720600.nc RapdD_al05.etrs.laea_19720700.nc RapdD_al05.etrs.laea_19720800.nc RapdD_al05.etrs.laea_19720900.nc RapdD_al05.etrs.laea_19721000.nc RapdD_al05.etrs.laea_19721100.nc RapdD_al05.etrs.laea_19721200.nc RapdD_al05.etrs.laea_19730100.nc RapdD_al05.etrs.laea_19730200.nc RapdD_al05.etrs.laea_19730300.nc RapdD_al05.etrs.laea_19730400.nc RapdD_al05.etrs.laea_19730500.nc RapdD_al05.etrs.laea_19730600.nc RapdD_al05.etrs.laea_19730700.nc RapdD_al05.etrs.laea_19730800.nc RapdD_al05.etrs.laea_19730900.nc RapdD_al05.etrs.laea_19731000.nc RapdD_al05.etrs.laea_19731100.nc RapdD_al05.etrs.laea_19731200.nc RapdD_al05.etrs.laea_19740100.nc RapdD_al05.etrs.laea_19740200.nc RapdD_al05.etrs.laea_19740300.nc RapdD_al05.etrs.laea_19740400.nc RapdD_al05.etrs.laea_19740500.nc RapdD_al05.etrs.laea_19740600.nc RapdD_al05.etrs.laea_19740700.nc RapdD_al05.etrs.laea_19740800.nc RapdD_al05.etrs.laea_19740900.nc RapdD_al05.etrs.laea_19741000.nc RapdD_al05.etrs.laea_19741100.nc RapdD_al05.etrs.laea_19741200.nc RapdD_al05.etrs.laea_19750100.nc RapdD_al05.etrs.laea_19750200.nc RapdD_al05.etrs.laea_19750300.nc RapdD_al05.etrs.laea_19750400.nc RapdD_al05.etrs.laea_19750500.nc RapdD_al05.etrs.laea_19750600.nc RapdD_al05.etrs.laea_19750700.nc RapdD_al05.etrs.laea_19750800.nc RapdD_al05.etrs.laea_19750900.nc RapdD_al05.etrs.laea_19751000.nc RapdD_al05.etrs.laea_19751100.nc RapdD_al05.etrs.laea_19751200.nc RapdD_al05.etrs.laea_19760100.nc RapdD_al05.etrs.laea_19760200.nc RapdD_al05.etrs.laea_19760300.nc RapdD_al05.etrs.laea_19760400.nc RapdD_al05.etrs.laea_19760500.nc RapdD_al05.etrs.laea_19760600.nc RapdD_al05.etrs.laea_19760700.nc RapdD_al05.etrs.laea_19760800.nc RapdD_al05.etrs.laea_19760900.nc RapdD_al05.etrs.laea_19761000.nc RapdD_al05.etrs.laea_19761100.nc RapdD_al05.etrs.laea_19761200.nc RapdD_al05.etrs.laea_19770100.nc RapdD_al05.etrs.laea_19770200.nc RapdD_al05.etrs.laea_19770300.nc RapdD_al05.etrs.laea_19770400.nc RapdD_al05.etrs.laea_19770500.nc RapdD_al05.etrs.laea_19770600.nc RapdD_al05.etrs.laea_19770700.nc RapdD_al05.etrs.laea_19770800.nc RapdD_al05.etrs.laea_19770900.nc RapdD_al05.etrs.laea_19771000.nc RapdD_al05.etrs.laea_19771100.nc RapdD_al05.etrs.laea_19771200.nc RapdD_al05.etrs.laea_19780100.nc RapdD_al05.etrs.laea_19780200.nc RapdD_al05.etrs.laea_19780300.nc RapdD_al05.etrs.laea_19780400.nc RapdD_al05.etrs.laea_19780500.nc RapdD_al05.etrs.laea_19780600.nc RapdD_al05.etrs.laea_19780700.nc RapdD_al05.etrs.laea_19780800.nc RapdD_al05.etrs.laea_19780900.nc RapdD_al05.etrs.laea_19781000.nc RapdD_al05.etrs.laea_19781100.nc RapdD_al05.etrs.laea_19781200.nc RapdD_al05.etrs.laea_19790100.nc RapdD_al05.etrs.laea_19790200.nc RapdD_al05.etrs.laea_19790300.nc RapdD_al05.etrs.laea_19790400.nc RapdD_al05.etrs.laea_19790500.nc RapdD_al05.etrs.laea_19790600.nc RapdD_al05.etrs.laea_19790700.nc RapdD_al05.etrs.laea_19790800.nc RapdD_al05.etrs.laea_19790900.nc RapdD_al05.etrs.laea_19791000.nc RapdD_al05.etrs.laea_19791100.nc RapdD_al05.etrs.laea_19791200.nc RapdD_al05.etrs.laea_19800100.nc RapdD_al05.etrs.laea_19800200.nc RapdD_al05.etrs.laea_19800300.nc RapdD_al05.etrs.laea_19800400.nc RapdD_al05.etrs.laea_19800500.nc RapdD_al05.etrs.laea_19800600.nc RapdD_al05.etrs.laea_19800700.nc RapdD_al05.etrs.laea_19800800.nc RapdD_al05.etrs.laea_19800900.nc RapdD_al05.etrs.laea_19801000.nc RapdD_al05.etrs.laea_19801100.nc RapdD_al05.etrs.laea_19801200.nc RapdD_al05.etrs.laea_19810100.nc RapdD_al05.etrs.laea_19810200.nc RapdD_al05.etrs.laea_19810300.nc RapdD_al05.etrs.laea_19810400.nc RapdD_al05.etrs.laea_19810500.nc RapdD_al05.etrs.laea_19810600.nc RapdD_al05.etrs.laea_19810700.nc RapdD_al05.etrs.laea_19810800.nc RapdD_al05.etrs.laea_19810900.nc RapdD_al05.etrs.laea_19811000.nc RapdD_al05.etrs.laea_19811100.nc RapdD_al05.etrs.laea_19811200.nc RapdD_al05.etrs.laea_19820100.nc RapdD_al05.etrs.laea_19820200.nc RapdD_al05.etrs.laea_19820300.nc RapdD_al05.etrs.laea_19820400.nc RapdD_al05.etrs.laea_19820500.nc RapdD_al05.etrs.laea_19820600.nc RapdD_al05.etrs.laea_19820700.nc RapdD_al05.etrs.laea_19820800.nc RapdD_al05.etrs.laea_19820900.nc RapdD_al05.etrs.laea_19821000.nc RapdD_al05.etrs.laea_19821100.nc RapdD_al05.etrs.laea_19821200.nc RapdD_al05.etrs.laea_19830100.nc RapdD_al05.etrs.laea_19830200.nc RapdD_al05.etrs.laea_19830300.nc RapdD_al05.etrs.laea_19830400.nc RapdD_al05.etrs.laea_19830500.nc RapdD_al05.etrs.laea_19830600.nc RapdD_al05.etrs.laea_19830700.nc RapdD_al05.etrs.laea_19830800.nc RapdD_al05.etrs.laea_19830900.nc RapdD_al05.etrs.laea_19831000.nc RapdD_al05.etrs.laea_19831100.nc RapdD_al05.etrs.laea_19831200.nc RapdD_al05.etrs.laea_19840100.nc RapdD_al05.etrs.laea_19840200.nc RapdD_al05.etrs.laea_19840300.nc RapdD_al05.etrs.laea_19840400.nc RapdD_al05.etrs.laea_19840500.nc RapdD_al05.etrs.laea_19840600.nc RapdD_al05.etrs.laea_19840700.nc RapdD_al05.etrs.laea_19840800.nc RapdD_al05.etrs.laea_19840900.nc RapdD_al05.etrs.laea_19841000.nc RapdD_al05.etrs.laea_19841100.nc RapdD_al05.etrs.laea_19841200.nc RapdD_al05.etrs.laea_19850100.nc RapdD_al05.etrs.laea_19850200.nc RapdD_al05.etrs.laea_19850300.nc RapdD_al05.etrs.laea_19850400.nc RapdD_al05.etrs.laea_19850500.nc RapdD_al05.etrs.laea_19850600.nc RapdD_al05.etrs.laea_19850700.nc RapdD_al05.etrs.laea_19850800.nc RapdD_al05.etrs.laea_19850900.nc RapdD_al05.etrs.laea_19851000.nc RapdD_al05.etrs.laea_19851100.nc RapdD_al05.etrs.laea_19851200.nc RapdD_al05.etrs.laea_19860100.nc RapdD_al05.etrs.laea_19860200.nc RapdD_al05.etrs.laea_19860300.nc RapdD_al05.etrs.laea_19860400.nc RapdD_al05.etrs.laea_19860500.nc RapdD_al05.etrs.laea_19860600.nc RapdD_al05.etrs.laea_19860700.nc RapdD_al05.etrs.laea_19860800.nc RapdD_al05.etrs.laea_19860900.nc RapdD_al05.etrs.laea_19861000.nc RapdD_al05.etrs.laea_19861100.nc RapdD_al05.etrs.laea_19861200.nc RapdD_al05.etrs.laea_19870100.nc RapdD_al05.etrs.laea_19870200.nc RapdD_al05.etrs.laea_19870300.nc RapdD_al05.etrs.laea_19870400.nc RapdD_al05.etrs.laea_19870500.nc RapdD_al05.etrs.laea_19870600.nc RapdD_al05.etrs.laea_19870700.nc RapdD_al05.etrs.laea_19870800.nc RapdD_al05.etrs.laea_19870900.nc RapdD_al05.etrs.laea_19871000.nc RapdD_al05.etrs.laea_19871100.nc RapdD_al05.etrs.laea_19871200.nc RapdD_al05.etrs.laea_19880100.nc RapdD_al05.etrs.laea_19880200.nc RapdD_al05.etrs.laea_19880300.nc RapdD_al05.etrs.laea_19880400.nc RapdD_al05.etrs.laea_19880500.nc RapdD_al05.etrs.laea_19880600.nc RapdD_al05.etrs.laea_19880700.nc RapdD_al05.etrs.laea_19880800.nc RapdD_al05.etrs.laea_19880900.nc RapdD_al05.etrs.laea_19881000.nc RapdD_al05.etrs.laea_19881100.nc RapdD_al05.etrs.laea_19881200.nc RapdD_al05.etrs.laea_19890100.nc RapdD_al05.etrs.laea_19890200.nc RapdD_al05.etrs.laea_19890300.nc RapdD_al05.etrs.laea_19890400.nc RapdD_al05.etrs.laea_19890500.nc RapdD_al05.etrs.laea_19890600.nc RapdD_al05.etrs.laea_19890700.nc RapdD_al05.etrs.laea_19890800.nc RapdD_al05.etrs.laea_19890900.nc RapdD_al05.etrs.laea_19891000.nc RapdD_al05.etrs.laea_19891100.nc RapdD_al05.etrs.laea_19891200.nc RapdD_al05.etrs.laea_19900100.nc RapdD_al05.etrs.laea_19900200.nc RapdD_al05.etrs.laea_19900300.nc RapdD_al05.etrs.laea_19900400.nc RapdD_al05.etrs.laea_19900500.nc RapdD_al05.etrs.laea_19900600.nc RapdD_al05.etrs.laea_19900700.nc RapdD_al05.etrs.laea_19900800.nc RapdD_al05.etrs.laea_19900900.nc RapdD_al05.etrs.laea_19901000.nc RapdD_al05.etrs.laea_19901100.nc RapdD_al05.etrs.laea_19901200.nc RapdD_al05.etrs.laea_19910100.nc RapdD_al05.etrs.laea_19910200.nc RapdD_al05.etrs.laea_19910300.nc RapdD_al05.etrs.laea_19910400.nc RapdD_al05.etrs.laea_19910500.nc RapdD_al05.etrs.laea_19910600.nc RapdD_al05.etrs.laea_19910700.nc RapdD_al05.etrs.laea_19910800.nc RapdD_al05.etrs.laea_19910900.nc RapdD_al05.etrs.laea_19911000.nc RapdD_al05.etrs.laea_19911100.nc RapdD_al05.etrs.laea_19911200.nc RapdD_al05.etrs.laea_19920100.nc RapdD_al05.etrs.laea_19920200.nc RapdD_al05.etrs.laea_19920300.nc RapdD_al05.etrs.laea_19920400.nc RapdD_al05.etrs.laea_19920500.nc RapdD_al05.etrs.laea_19920600.nc RapdD_al05.etrs.laea_19920700.nc RapdD_al05.etrs.laea_19920800.nc RapdD_al05.etrs.laea_19920900.nc RapdD_al05.etrs.laea_19921000.nc RapdD_al05.etrs.laea_19921100.nc RapdD_al05.etrs.laea_19921200.nc RapdD_al05.etrs.laea_19930100.nc RapdD_al05.etrs.laea_19930200.nc RapdD_al05.etrs.laea_19930300.nc RapdD_al05.etrs.laea_19930400.nc RapdD_al05.etrs.laea_19930500.nc RapdD_al05.etrs.laea_19930600.nc RapdD_al05.etrs.laea_19930700.nc RapdD_al05.etrs.laea_19930800.nc RapdD_al05.etrs.laea_19930900.nc RapdD_al05.etrs.laea_19931000.nc RapdD_al05.etrs.laea_19931100.nc RapdD_al05.etrs.laea_19931200.nc RapdD_al05.etrs.laea_19940100.nc RapdD_al05.etrs.laea_19940200.nc RapdD_al05.etrs.laea_19940300.nc RapdD_al05.etrs.laea_19940400.nc RapdD_al05.etrs.laea_19940500.nc RapdD_al05.etrs.laea_19940600.nc RapdD_al05.etrs.laea_19940700.nc RapdD_al05.etrs.laea_19940800.nc RapdD_al05.etrs.laea_19940900.nc RapdD_al05.etrs.laea_19941000.nc RapdD_al05.etrs.laea_19941100.nc RapdD_al05.etrs.laea_19941200.nc RapdD_al05.etrs.laea_19950100.nc RapdD_al05.etrs.laea_19950200.nc RapdD_al05.etrs.laea_19950300.nc RapdD_al05.etrs.laea_19950400.nc RapdD_al05.etrs.laea_19950500.nc RapdD_al05.etrs.laea_19950600.nc RapdD_al05.etrs.laea_19950700.nc RapdD_al05.etrs.laea_19950800.nc RapdD_al05.etrs.laea_19950900.nc RapdD_al05.etrs.laea_19951000.nc RapdD_al05.etrs.laea_19951100.nc RapdD_al05.etrs.laea_19951200.nc RapdD_al05.etrs.laea_19960100.nc RapdD_al05.etrs.laea_19960200.nc RapdD_al05.etrs.laea_19960300.nc RapdD_al05.etrs.laea_19960400.nc RapdD_al05.etrs.laea_19960500.nc RapdD_al05.etrs.laea_19960600.nc RapdD_al05.etrs.laea_19960700.nc RapdD_al05.etrs.laea_19960800.nc RapdD_al05.etrs.laea_19960900.nc RapdD_al05.etrs.laea_19961000.nc RapdD_al05.etrs.laea_19961100.nc RapdD_al05.etrs.laea_19961200.nc RapdD_al05.etrs.laea_19970100.nc RapdD_al05.etrs.laea_19970200.nc RapdD_al05.etrs.laea_19970300.nc RapdD_al05.etrs.laea_19970400.nc RapdD_al05.etrs.laea_19970500.nc RapdD_al05.etrs.laea_19970600.nc RapdD_al05.etrs.laea_19970700.nc RapdD_al05.etrs.laea_19970800.nc RapdD_al05.etrs.laea_19970900.nc RapdD_al05.etrs.laea_19971000.nc RapdD_al05.etrs.laea_19971100.nc RapdD_al05.etrs.laea_19971200.nc RapdD_al05.etrs.laea_19980100.nc RapdD_al05.etrs.laea_19980200.nc RapdD_al05.etrs.laea_19980300.nc RapdD_al05.etrs.laea_19980400.nc RapdD_al05.etrs.laea_19980500.nc RapdD_al05.etrs.laea_19980600.nc RapdD_al05.etrs.laea_19980700.nc RapdD_al05.etrs.laea_19980800.nc RapdD_al05.etrs.laea_19980900.nc RapdD_al05.etrs.laea_19981000.nc RapdD_al05.etrs.laea_19981100.nc RapdD_al05.etrs.laea_19981200.nc RapdD_al05.etrs.laea_19990100.nc RapdD_al05.etrs.laea_19990200.nc RapdD_al05.etrs.laea_19990300.nc RapdD_al05.etrs.laea_19990400.nc RapdD_al05.etrs.laea_19990500.nc RapdD_al05.etrs.laea_19990600.nc RapdD_al05.etrs.laea_19990700.nc RapdD_al05.etrs.laea_19990800.nc RapdD_al05.etrs.laea_19990900.nc RapdD_al05.etrs.laea_19991000.nc RapdD_al05.etrs.laea_19991100.nc RapdD_al05.etrs.laea_19991200.nc RapdD_al05.etrs.laea_20000100.nc RapdD_al05.etrs.laea_20000200.nc RapdD_al05.etrs.laea_20000300.nc RapdD_al05.etrs.laea_20000400.nc RapdD_al05.etrs.laea_20000500.nc RapdD_al05.etrs.laea_20000600.nc RapdD_al05.etrs.laea_20000700.nc RapdD_al05.etrs.laea_20000800.nc RapdD_al05.etrs.laea_20000900.nc RapdD_al05.etrs.laea_20001000.nc RapdD_al05.etrs.laea_20001100.nc RapdD_al05.etrs.laea_20001200.nc RapdD_al05.etrs.laea_20010100.nc RapdD_al05.etrs.laea_20010200.nc RapdD_al05.etrs.laea_20010300.nc RapdD_al05.etrs.laea_20010400.nc RapdD_al05.etrs.laea_20010500.nc RapdD_al05.etrs.laea_20010600.nc RapdD_al05.etrs.laea_20010700.nc RapdD_al05.etrs.laea_20010800.nc RapdD_al05.etrs.laea_20010900.nc RapdD_al05.etrs.laea_20011000.nc RapdD_al05.etrs.laea_20011100.nc RapdD_al05.etrs.laea_20011200.nc RapdD_al05.etrs.laea_20020100.nc RapdD_al05.etrs.laea_20020200.nc RapdD_al05.etrs.laea_20020300.nc RapdD_al05.etrs.laea_20020400.nc RapdD_al05.etrs.laea_20020500.nc RapdD_al05.etrs.laea_20020600.nc RapdD_al05.etrs.laea_20020700.nc RapdD_al05.etrs.laea_20020800.nc RapdD_al05.etrs.laea_20020900.nc RapdD_al05.etrs.laea_20021000.nc RapdD_al05.etrs.laea_20021100.nc RapdD_al05.etrs.laea_20021200.nc RapdD_al05.etrs.laea_20030100.nc RapdD_al05.etrs.laea_20030200.nc RapdD_al05.etrs.laea_20030300.nc RapdD_al05.etrs.laea_20030400.nc RapdD_al05.etrs.laea_20030500.nc RapdD_al05.etrs.laea_20030600.nc RapdD_al05.etrs.laea_20030700.nc RapdD_al05.etrs.laea_20030800.nc RapdD_al05.etrs.laea_20030900.nc RapdD_al05.etrs.laea_20031000.nc RapdD_al05.etrs.laea_20031100.nc RapdD_al05.etrs.laea_20031200.nc RapdD_al05.etrs.laea_20040100.nc RapdD_al05.etrs.laea_20040200.nc RapdD_al05.etrs.laea_20040300.nc RapdD_al05.etrs.laea_20040400.nc RapdD_al05.etrs.laea_20040500.nc RapdD_al05.etrs.laea_20040600.nc RapdD_al05.etrs.laea_20040700.nc RapdD_al05.etrs.laea_20040800.nc RapdD_al05.etrs.laea_20040900.nc RapdD_al05.etrs.laea_20041000.nc RapdD_al05.etrs.laea_20041100.nc RapdD_al05.etrs.laea_20041200.nc RapdD_al05.etrs.laea_20050100.nc RapdD_al05.etrs.laea_20050200.nc RapdD_al05.etrs.laea_20050300.nc RapdD_al05.etrs.laea_20050400.nc RapdD_al05.etrs.laea_20050500.nc RapdD_al05.etrs.laea_20050600.nc RapdD_al05.etrs.laea_20050700.nc RapdD_al05.etrs.laea_20050800.nc RapdD_al05.etrs.laea_20050900.nc RapdD_al05.etrs.laea_20051000.nc RapdD_al05.etrs.laea_20051100.nc RapdD_al05.etrs.laea_20051200.nc RapdD_al05.etrs.laea_20060100.nc RapdD_al05.etrs.laea_20060200.nc RapdD_al05.etrs.laea_20060300.nc RapdD_al05.etrs.laea_20060400.nc RapdD_al05.etrs.laea_20060500.nc RapdD_al05.etrs.laea_20060600.nc RapdD_al05.etrs.laea_20060700.nc RapdD_al05.etrs.laea_20060800.nc RapdD_al05.etrs.laea_20060900.nc RapdD_al05.etrs.laea_20061000.nc RapdD_al05.etrs.laea_20061100.nc RapdD_al05.etrs.laea_20061200.nc RapdD_al05.etrs.laea_20070100.nc RapdD_al05.etrs.laea_20070200.nc RapdD_al05.etrs.laea_20070300.nc RapdD_al05.etrs.laea_20070400.nc RapdD_al05.etrs.laea_20070500.nc RapdD_al05.etrs.laea_20070600.nc RapdD_al05.etrs.laea_20070700.nc RapdD_al05.etrs.laea_20070800.nc RapdD_al05.etrs.laea_20070900.nc RapdD_al05.etrs.laea_20071000.nc RapdD_al05.etrs.laea_20071100.nc RapdD_al05.etrs.laea_20071200.nc RapdD_al05.etrs.laea_20080100.nc RapdD_al05.etrs.laea_20080200.nc RapdD_al05.etrs.laea_20080300.nc RapdD_al05.etrs.laea_20080400.nc RapdD_al05.etrs.laea_20080500.nc RapdD_al05.etrs.laea_20080600.nc RapdD_al05.etrs.laea_20080700.nc RapdD_al05.etrs.laea_20080800.nc RapdD_al05.etrs.laea_20080900.nc RapdD_al05.etrs.laea_20081000.nc RapdD_al05.etrs.laea_20081100.nc RapdD_al05.etrs.laea_20081200.nc EURO4M-APGD-1971-2008.nc" ;
		:institution = "Federal Office of Meteorology and Climatology MeteoSwiss" ;
		:Conventions = "CF-1.4" ;
		:References = "Isotta, F.A. et al. 2013: The climate of daily precipitation in the Alps: development and analysis of a high-resolution grid dataset from pan-Alpine rain-gauge data. Int. J. Climatol., accepted. Please check for updates on the publication status!" ;
		:nco_openmp_thread_number = 1 ;
		:CDO = "Climate Data Operators version 1.9.1 (http://mpimet.mpg.de/cdo)" ;
}
